netcdf roms_frc {
dimensions:
	xi_rho = 12 ;
	xi_u = 11 ;
	xi_v = 12 ;
	xi_psi = 11 ;
	eta_rho = 14 ;
	eta_u = 14 ;
	eta_v = 13 ;
	eta_psi = 13 ;
	ocean_time = 2 ; // (2 currently)
variables:
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 1970-01-01 00:00:00" ;
		ocean_time:calendar = "proleptic_gregorian" ;
		ocean_time:field = "time, scalar, series" ;
	float shflux(ocean_time, eta_rho, xi_rho) ;
		shflux:long_name = "surface net heat flux" ;
		shflux:units = "watt meter-2" ;
		shflux:negative_value = "upward flux, cooling" ;
		shflux:positive_value = "downward flux, heating" ;
		shflux:time = "ocean_time" ;
		shflux:grid = "grid" ;
		shflux:location = "face" ;
		shflux:coordinates = "x_rho y_rho ocean_time" ;
		shflux:field = "surface heat flux, scalar, series" ;
	float swflux(ocean_time, eta_rho, xi_rho) ;
		swflux:long_name = "surface net freshwater flux, (E-P)" ;
		swflux:units = "meter second-1" ;
		swflux:time = "ocean_time" ;
		swflux:grid = "grid" ;
		swflux:location = "face" ;
		swflux:coordinates = "x_rho y_rho ocean_time" ;
		swflux:field = "surface net freshwater flux, scalar, series" ;
	float swrad(ocean_time, eta_rho, xi_rho) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:negative_value = "upward flux, cooling" ;
		swrad:positive_value = "downward flux, heating" ;
		swrad:time = "ocean_time" ;
		swrad:grid = "grid" ;
		swrad:location = "face" ;
		swrad:coordinates = "x_rho y_rho ocean_time" ;
		swrad:field = "shortwave radiation, scalar, series" ;
	float sustr(ocean_time, eta_u, xi_u) ;
		sustr:long_name = "surface u-momentum stress" ;
		sustr:units = "newton meter-2" ;
		sustr:time = "ocean_time" ;
		sustr:grid = "grid" ;
		sustr:location = "edge1" ;
		sustr:coordinates = "x_u y_u ocean_time" ;
		sustr:field = "surface u-momentum stress, scalar, series" ;
	float svstr(ocean_time, eta_v, xi_v) ;
		svstr:long_name = "surface v-momentum stress" ;
		svstr:units = "newton meter-2" ;
		svstr:time = "ocean_time" ;
		svstr:grid = "grid" ;
		svstr:location = "edge2" ;
		svstr:coordinates = "x_v y_v ocean_time" ;
		svstr:field = "surface v-momentum stress, scalar, series" ;

// global attributes:
		:file = "roms_frc.nc" ;
		:format = "netCDF-3 64bit offset file" ;
		:Conventions = "CF-1.4, SGRID-0.3" ;
		:type = "ROMS/TOMS history file" ;
		:title = "Column model for turbulence scheme testing" ;
		:var_info = "../External/varinfo.dat" ;
		:svn_url = "https://www.myroms.org/svn/src/trunk" ;
		:svn_rev = "986" ;
		:code_dir = "/home/kaihc/ROMS-trunk" ;
		:header_dir = "/home/kaihc/Desktop/R1D/Include" ;
		:header_file = "column.h" ;
		:os = "Linux" ;
		:cpu = "x86_64" ;
		:compiler_system = "gfortran" ;
		:compiler_command = "/usr/bin/gfortran" ;
		:compiler_flags = "-frepack-arrays -O3 -ffast-math -" ;
}
