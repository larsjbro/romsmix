netcdf ocean_frc_800m_2018 {
dimensions:
	ocean_time = UNLIMITED ; // (2920 currently)
	eta_rho = 1148 ;
	xi_rho = 2747 ;
variables:
	float rain(ocean_time, eta_rho, xi_rho) ;
		rain:coordinates = "lon lat" ;
		rain:grid_mapping = "projection_stere" ;
		rain:standard_name = "lwe_thickness_of_percipitation_amount" ;
		rain:units = "kg/m2/s" ;
		rain:cell_methods = "surface: mean" ;
	double Qair(ocean_time, eta_rho, xi_rho) ;
		Qair:coordinates = "lon lat" ;
		Qair:grid_mapping = "projection_stere" ;
		Qair:units = "percentage" ;
		Qair:cell_methods = "surface: mean" ;
	float dewpoint(ocean_time, eta_rho, xi_rho) ;
		dewpoint:coordinates = "lon lat" ;
		dewpoint:grid_mapping = "projection_stere" ;
		dewpoint:units = "C" ;
		dewpoint:cell_methods = "surface: mean" ;
	float Tair(ocean_time, eta_rho, xi_rho) ;
		Tair:coordinates = "lon lat" ;
		Tair:grid_mapping = "projection_stere" ;
		Tair:standard_name = "air_temperature" ;
		Tair:units = "C" ;
		Tair:cell_methods = "surface: mean" ;
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "time" ;
		ocean_time:standard_name = "time" ;
		ocean_time:units = "days since 1970-01-01 00:00:00 +00:00" ;
	double forecast_reference_time ;
		forecast_reference_time:units = "seconds since 1970-01-01 00:00:00 +00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
	short surface ;
		surface:_FillValue = -32767s ;
		surface:description = "ground or water surface" ;
		surface:long_name = "surface" ;
		surface:positive = "up" ;
		surface:units = "m" ;
		surface:cell_methods = "surface: mean" ;
	float Pair(ocean_time, eta_rho, xi_rho) ;
		Pair:standard_name = "air_pressure_at_sea_level" ;
		Pair:units = "hPa" ;
		Pair:coordinates = "lon lat" ;
		Pair:grid_mapping = "projection_stere" ;
		Pair:cell_methods = "surface: mean" ;
	float cloud(ocean_time, eta_rho, xi_rho) ;
		cloud:standard_name = "cloud_area_fraction" ;
		cloud:units = "1" ;
		cloud:coordinates = "lon lat" ;
		cloud:grid_mapping = "projection_stere" ;
		cloud:cell_methods = "surface: mean" ;
	float Uwind(ocean_time, eta_rho, xi_rho) ;
		Uwind:standard_name = "x_wind" ;
		Uwind:units = "m/s" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:grid_mapping = "projection_stere" ;
		Uwind:cell_methods = "surface: mean" ;
	float Vwind(ocean_time, eta_rho, xi_rho) ;
		Vwind:standard_name = "y_wind" ;
		Vwind:units = "m/s" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:grid_mapping = "projection_stere" ;
		Vwind:cell_methods = "surface: mean" ;
	int projection_stere ;
		projection_stere:grid_mapping_name = "polar_stereographic" ;
		projection_stere:scale_factor_at_projection_origin = 0.933012701892219 ;
		projection_stere:straight_vertical_longitude_from_pole = 70. ;
		projection_stere:latitude_of_projection_origin = 90. ;
		projection_stere:false_easting = 3371200. ;
		projection_stere:false_northing = 1846400. ;
		projection_stere:semi_major_axis = 6378137. ;
		projection_stere:semi_minor_axis = 6356752.3142 ;
		projection_stere:proj4 = "+proj=stere +ellps=WGS84 +lat_0=90.0 +lat_ts=60.0 +x_0=3371200 +y_0=1846400 +lon_0=70" ;
	double xi_rho(xi_rho) ;
		xi_rho:standard_name = "projection_x_coordinate" ;
		xi_rho:units = "m" ;
	double eta_rho(eta_rho) ;
		eta_rho:standard_name = "projection_y_coordinate" ;
		eta_rho:units = "m" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:units = "degree_east" ;
		lon_rho:long_name = "longitude" ;
		lon_rho:standard_name = "longitude" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:units = "degree_north" ;
		lat_rho:long_name = "latitude" ;
		lat_rho:standard_name = "latitude" ;

// global attributes:
		:institution = "Norwegian Meteorological Institute, met.no" ;
		:source = "HIRLAM" ;
		:min_time = "2018-01-01 03:00:00Z" ;
		:max_time = "2018-01-01" ;
		:email = "kaihc@met.no" ;
		:history = "Sun Oct 11 21:00:29 2020: ncrcat /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_001.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_002.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_003.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_004.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_005.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_006.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_007.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_008.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_009.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_010.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_011.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_012.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_013.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_014.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_015.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_016.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_017.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_018.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_019.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_020.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_021.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_022.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_023.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_024.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_025.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_026.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_027.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_028.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_029.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_030.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_031.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_032.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_033.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_034.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_035.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_036.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_037.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_038.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_039.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_040.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_041.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_042.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_043.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_044.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_045.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_046.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_047.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_048.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_049.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_050.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_051.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_052.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_053.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_054.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_055.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_056.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_057.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_058.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_059.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_060.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_061.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_062.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_063.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_064.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_065.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_066.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_067.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_068.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_069.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_070.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_071.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_072.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_073.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_074.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_075.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_076.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_077.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_078.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_079.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_080.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_081.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_082.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_083.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_084.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_085.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_086.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_087.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_088.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_089.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_090.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_091.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_092.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_093.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_094.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_095.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_096.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_097.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_098.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_099.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_100.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_101.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_102.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_103.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_104.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_105.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_106.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_107.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_108.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_109.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_110.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_111.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_112.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_113.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_114.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_115.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_116.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_117.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_118.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_119.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_120.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_121.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_122.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_123.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_124.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_125.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_126.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_127.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_128.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_129.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_130.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_131.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_132.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_133.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_134.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_135.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_136.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_137.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_138.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_139.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_140.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_141.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_142.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_143.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_144.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_145.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_146.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_147.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_148.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_149.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_150.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_151.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_152.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_153.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_154.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_155.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_156.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_157.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_158.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_159.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_160.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_161.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_162.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_163.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_164.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_165.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_166.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_167.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_168.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_169.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_170.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_171.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_172.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_173.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_174.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_175.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_176.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_177.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_178.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_179.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_180.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_181.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_182.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_183.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_184.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_185.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_186.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_187.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_188.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_189.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_190.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_191.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_192.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_193.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_194.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_195.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_196.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_197.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_198.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_199.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_200.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_201.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_202.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_203.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_204.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_205.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_206.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_207.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_208.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_209.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_210.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_211.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_212.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_213.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_214.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_215.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_216.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_217.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_218.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_219.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_220.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_221.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_222.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_223.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_224.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_225.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_226.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_227.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_228.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_229.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_230.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_231.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_232.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_233.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_234.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_235.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_236.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_237.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_238.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_239.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_240.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_241.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_242.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_243.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_244.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_245.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_246.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_247.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_248.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_249.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_250.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_251.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_252.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_253.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_254.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_255.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_256.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_257.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_258.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_259.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_260.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_261.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_262.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_263.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_264.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_265.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_266.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_267.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_268.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_269.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_270.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_271.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_272.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_273.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_274.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_275.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_276.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_277.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_278.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_279.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_280.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_281.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_282.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_283.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_284.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_285.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_286.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_287.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_288.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_289.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_290.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_291.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_292.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_293.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_294.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_295.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_296.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_297.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_298.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_299.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_300.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_301.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_302.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_303.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_304.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_305.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_306.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_307.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_308.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_309.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_310.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_311.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_312.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_313.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_314.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_315.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_316.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_317.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_318.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_319.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_320.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_321.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_322.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_323.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_324.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_325.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_326.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_327.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_328.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_329.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_330.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_331.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_332.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_333.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_334.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_335.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_336.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_337.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_338.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_339.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_340.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_341.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_342.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_343.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_344.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_345.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_346.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_347.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_348.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_349.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_350.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_351.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_352.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_353.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_354.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_355.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_356.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_357.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_358.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_359.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_360.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_361.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_362.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_363.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_364.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_365.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/ocean_frc_800m_2018.nc\n",
			"Thu Oct  8 12:03:13 2020: ncrcat -O /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/forecast_00_001.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/forecast_12_001.nc -o /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/daily_001.nc\n",
			"Thu Oct  8 12:02:00 2020: ncrename -d latitude,eta_rho -d longitude,xi_rho /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/forecast_00_001.nc\n",
			"Thu Oct  8 12:01:56 2020: ncrename -v lat,lat_rho -v lon,lon_rho -v longitude,xi_rho -v latitude,eta_rho /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/forecast_00_001.nc\n",
			"Thu Oct  8 12:01:48 2020: ncwa -O -a surface /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/tmp.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/forecast_00_001.nc\n",
			"Thu Oct  8 12:01:34 2020: ncatted -a units,Qair,m,c,percentage /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/tmp.nc\n",
			"Thu Oct  8 12:01:25 2020: ncap2 -O -s Qair = 100*exp(17.502*( (dewpoint/(240.97+dewpoint)) - (Tair/(240.97+Tair)) )) /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/tmp.nc /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/tmp.nc\n",
			"Thu Oct  8 12:01:24 2020: ncatted -a units,Tair,m,c,C -a units,dewpoint,m,c,C /lustre/storeB/project/fou/hi/roms_operational/norkyst_v3/norkyst_DA/Forcing/tmp.nc\n",
			"2020-10-08 creation by fimex" ;
		:Conventions = "CF-1.0" ;
		:NCO = "\"4.5.4\"" ;
		:nco_openmp_thread_number = 1 ;
}
